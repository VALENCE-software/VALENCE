  1 1   1 0 1  12 4 1   5 21 0   0 0 0   1

  20 20 20   0 0 0  0.0 0.0



  1   0.0    0.0   0.0



  4.0   5
0   9
    14630.0000000              0.0000920        
     2191.0000000              0.0007130        
      498.2000000              0.0037350        
      140.9000000              0.0154680        
       45.8600000              0.0528740        
       16.4700000              0.1456940        
        6.3190000              0.3026810        
        2.5350000              0.4049360        
        1.0350000              0.2223870        
0   9
    14630.0000000             -0.0000170        
     2191.0000000             -0.0001300        
      498.2000000             -0.0006790        
      140.9000000             -0.0028570        
       45.8600000             -0.0098130        
       16.4700000             -0.0286090        
        6.3190000             -0.0637600        
        2.5350000             -0.1172310        
        1.0350000             -0.1212020        
0   1
        0.2528000                     
0   1
        0.1052000                     
0   1
        0.0426100                     


 1 2


      1        1   4
   2   -0.41969734   3   -0.65789598   4   -0.40843774   5   -0.10162906
      1        1   4
   2   -0.16546626   3    0.15183593   4   -0.68009037   5   -0.49468748
      1        1   4
   1    0.99439744   2    0.00032620   3    0.01226384   4    0.00233721


Beryllium atom ground state, 1s1s2s2s' singlet-S.
The above input is the same as the 'be' example except that the valence, 2s, orbital is 'split' into a spin-coupled pair, denoted 2s2s', and the wave function has been re-optimized.
(the above orbitals are optimized to 1d-6 kCal/Mol in the total energy, output given below)

 guess energy in atomic units          -14.5763526671383907

The energy is lower than the VSHF energy, reflecting a static correlation in the single-reference wave function.

